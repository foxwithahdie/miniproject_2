module top #(
    parameter c_PWM_INTERVAL = 1200
)(
    input logic clk,
    output logic RGB_R,
    output logic RGB_G,
    output logic RGB_B
);

initial begin

end

endmodule
`timescale 10ns/10ns
`include "../src/top.sv"

module test_top;

endmodule